`timescale 1ns/1ns
module vga_pic(
  input  wire        vga_clk,
  input  wire        sys_rst_n,
  input  wire [9:0]  pix_x,
  input  wire [9:0]  pix_y,
  output reg  [15:0] pix_data
);
  parameter   CHAR_B_H = 10'd140,
              CHAR_B_V = 10'd216,
              CHAR_W   = 10'd256,
              CHAR_H   = 10'd64,
              BLACK    = 16'h0000,
              WHITE    = 16'hFFFF,
              GOLDEN   = 16'hFEC0,
              PINK     = 16'hEE38;

  localparam integer BYTES_PER_ROW = CHAR_W/8;
  localparam integer ROM_SIZE      = CHAR_H*BYTES_PER_ROW;
  
    localparam [ROM_SIZE*8-1:0] ROMBITS = {
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b11111111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b01111111, 8'b11100000, 8'b00000000, 8'b00001111, 8'b11111100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111111, 8'b11111111, 8'b10000011, 8'b11111111, 8'b11111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011111, 8'b11111111, 8'b11101111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b01111111, 8'b11100000, 8'b00000000, 8'b00001111, 8'b11111100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111111, 8'b11111111, 8'b10000011, 8'b11111111, 8'b11111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111111, 8'b11111111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b01111111, 8'b11110000, 8'b00000000, 8'b00011111, 8'b11111100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111111, 8'b11111111, 8'b10000011, 8'b11111111, 8'b11111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111111, 8'b11001111, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b11111111, 8'b11111111, 8'b11111111, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11110000, 8'b00000000, 8'b00011111, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111110, 8'b00000000, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b00000000, 8'b01111000, 8'b00000011, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11110000, 8'b00000000, 8'b00111111, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b11111000, 8'b00000000, 8'b01111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b00000000, 8'b01111000, 8'b00000011, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11111000, 8'b00000000, 8'b00111111, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b11110000, 8'b00000000, 8'b00111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b00000000, 8'b01111000, 8'b00000011, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11111000, 8'b00000000, 8'b00111101, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b11100000, 8'b00000000, 8'b00011111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b00000000, 8'b01111000, 8'b00000011, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b01111100, 8'b00000000, 8'b01111101, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b11100000, 8'b00000000, 8'b00011111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b00000000, 8'b01111000, 8'b00000011, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b01111100, 8'b00000000, 8'b01111101, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11100000, 8'b00000000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b00000000, 8'b01111000, 8'b00000011, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00111110, 8'b00000000, 8'b11111001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11100000, 8'b00000000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b00000000, 8'b01111000, 8'b00000011, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00111110, 8'b00000000, 8'b11111001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11100000, 8'b00000000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b00000000, 8'b01111000, 8'b00000011, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00011111, 8'b00000001, 8'b11110001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b00000000, 8'b01111000, 8'b00000011, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00011111, 8'b00000001, 8'b11110001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b00000000, 8'b01111000, 8'b00000001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00001111, 8'b00000001, 8'b11100001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b11111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b00000000, 8'b01111000, 8'b00000001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00001111, 8'b10000011, 8'b11100001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00001111, 8'b10000011, 8'b11100001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111111, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00000111, 8'b11000111, 8'b11000001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111111, 8'b11111111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00000111, 8'b11000111, 8'b11000001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b11111111, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00000011, 8'b11101111, 8'b10000001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b11111111, 8'b11111100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00000011, 8'b11101111, 8'b10000001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011111, 8'b11111110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00000001, 8'b11101111, 8'b00000001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00000001, 8'b11111111, 8'b00000001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00000000, 8'b11111111, 8'b00000001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00000000, 8'b11111110, 8'b00000001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00000000, 8'b11111110, 8'b00000001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00000000, 8'b01111100, 8'b00000001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00001111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00000000, 8'b00000000, 8'b00000001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11100000, 8'b00000000, 8'b00001111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00000000, 8'b00000000, 8'b00000001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11100000, 8'b00000000, 8'b00001111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00000000, 8'b00000000, 8'b00000001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11100000, 8'b00000000, 8'b00011111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00000000, 8'b00000000, 8'b00000001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b11110000, 8'b00000000, 8'b00011111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b11100000, 8'b00000000, 8'b00001111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00000000, 8'b00000000, 8'b00000001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b11111000, 8'b00000000, 8'b00111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b11110000, 8'b00000000, 8'b00001111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00000000, 8'b00000000, 8'b00000001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111100, 8'b00000000, 8'b01111110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b11111000, 8'b00000000, 8'b00111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b00000000, 8'b00000000, 8'b00000001, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111110, 8'b00000001, 8'b11111100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b11111100, 8'b00000000, 8'b01111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b11111111, 8'b11111110, 8'b00000000, 8'b11111111, 8'b11111110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111111, 8'b11001111, 8'b11111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b11111111, 8'b11000111, 8'b11111110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111111, 8'b11111111, 8'b11111100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b11111111, 8'b11111110, 8'b00000000, 8'b11111111, 8'b11111110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111111, 8'b11111111, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b10111111, 8'b11111111, 8'b11111100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111111, 8'b11111111, 8'b11111100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b11111111, 8'b11111110, 8'b00000000, 8'b11111111, 8'b11111110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b11111111, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b10011111, 8'b11111111, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111111, 8'b11111111, 8'b11111100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11111111, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b11111111, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
};
  reg [7:0] bmp [0:ROM_SIZE-1];

  integer i;
  reg [ROM_SIZE*8-1:0] tmp;
  initial begin
    tmp = ROMBITS;
    for (i = 0; i < ROM_SIZE; i = i + 1) begin
      bmp[i] = tmp[ROM_SIZE*8-1 : ROM_SIZE*8-8];
      tmp    = {tmp[ROM_SIZE*8-9:0], 8'b00000000};
    end
  end

  wire in_box;
  wire [9:0] x, y;
  wire [10:0] byte_idx;
  wire [2:0]  bit_idx;
  wire        bit_on;

  assign in_box  = (pix_x >= CHAR_B_H) && (pix_x < CHAR_B_H + CHAR_W) &&
                   (pix_y >= CHAR_B_V) && (pix_y < CHAR_B_V + CHAR_H);
  assign x = pix_x - CHAR_B_H;
  assign y = pix_y - CHAR_B_V;

  assign byte_idx = y*BYTES_PER_ROW + (x >> 3);
  assign bit_idx  = 3'd7 - x[2:0];
  assign bit_on   = bmp[byte_idx][bit_idx];

  always @(posedge vga_clk or negedge sys_rst_n) begin
    if(!sys_rst_n)             pix_data <= BLACK;
    else if(in_box && bit_on)  pix_data <= PINK;
    else                       pix_data <= BLACK;
  end
endmodule