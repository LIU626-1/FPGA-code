`timescale 1ns/1ns
module tb_Running_light();

reg sys_clk;
reg sys_rst_n;
wire led0;
wire led1;
wire led2;
wire led3;

initial begin
 sys_clk = 1'b1;
 sys_rst_n <= 1'b0;
 #20
 sys_rst_n <= 1'b1;
end

always #10 sys_clk = ~sys_clk;

Running_light Running_light_instance(
 .sys_clk (sys_clk),
 .sys_rst_n (sys_rst_n),
 .led0(led0),
 .led1(led1),
 .led2(led2),
 .led3(led3)
);

endmodule